module top(input [3:0] bus);
endmodule //top
